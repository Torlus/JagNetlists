/* verilator lint_off LITENDIAN */
`include "defs.v"

module j_jbus
(
	input ain_0,
	input ain_1,
	input ain_2,
	input ain_3,
	input ain_4,
	input ain_5,
	input ain_6,
	input ain_7,
	input ain_8,
	input ain_9,
	input ain_10,
	input ain_11,
	input ain_12,
	input ain_13,
	input ain_14,
	input ain_15,
	input ain_16,
	input ain_17,
	input ain_18,
	input ain_19,
	input ain_20,
	input ain_21,
	input ain_22,
	input ain_23,
	input din_0,
	input din_1,
	input din_2,
	input din_3,
	input din_4,
	input din_5,
	input din_6,
	input din_7,
	input din_8,
	input din_9,
	input din_10,
	input din_11,
	input din_12,
	input din_13,
	input din_14,
	input din_15,
	input din_16,
	input din_17,
	input din_18,
	input din_19,
	input din_20,
	input din_21,
	input din_22,
	input din_23,
	input din_24,
	input din_25,
	input din_26,
	input din_27,
	input din_28,
	input din_29,
	input din_30,
	input din_31,
	input dr_0,
	input dr_1,
	input dr_2,
	input dr_3,
	input dr_4,
	input dr_5,
	input dr_6,
	input dr_7,
	input dr_8,
	input dr_9,
	input dr_10,
	input dr_11,
	input dr_12,
	input dr_13,
	input dr_14,
	input dr_15,
	input dinlatch_0,
	input dinlatch_1,
	input dmuxd_0,
	input dmuxd_1,
	input dmuxu_0,
	input dmuxu_1,
	input dren,
	input xdsrc,
	input ack,
	input wd_0,
	input wd_1,
	input wd_2,
	input wd_3,
	input wd_4,
	input wd_5,
	input wd_6,
	input wd_7,
	input wd_8,
	input wd_9,
	input wd_10,
	input wd_11,
	input wd_12,
	input wd_13,
	input wd_14,
	input wd_15,
	input wd_16,
	input wd_17,
	input wd_18,
	input wd_19,
	input wd_20,
	input wd_21,
	input wd_22,
	input wd_23,
	input wd_24,
	input wd_25,
	input wd_26,
	input wd_27,
	input wd_28,
	input wd_29,
	input wd_30,
	input wd_31,
	input clk,
	input cfg_0,
	input cfg_1,
	input cfgw,
	input a_0,
	input a_1,
	input a_2,
	input a_3,
	input a_4,
	input a_5,
	input a_6,
	input a_7,
	input a_8,
	input a_9,
	input a_10,
	input a_11,
	input a_12,
	input a_13,
	input a_14,
	input a_15,
	input a_16,
	input a_17,
	input a_18,
	input a_19,
	input a_20,
	input a_21,
	input a_22,
	input a_23,
	input ainen,
	input seta1,
	input masterdata,
	output dout_0,
	output dout_1,
	output dout_2,
	output dout_3,
	output dout_4,
	output dout_5,
	output dout_6,
	output dout_7,
	output dout_8,
	output dout_9,
	output dout_10,
	output dout_11,
	output dout_12,
	output dout_13,
	output dout_14,
	output dout_15,
	output dout_16,
	output dout_17,
	output dout_18,
	output dout_19,
	output dout_20,
	output dout_21,
	output dout_22,
	output dout_23,
	output dout_24,
	output dout_25,
	output dout_26,
	output dout_27,
	output dout_28,
	output dout_29,
	output dout_30,
	output dout_31,
	output aout_0,
	output aout_1,
	output aout_2,
	output aout_3,
	output aout_4,
	output aout_5,
	output aout_6,
	output aout_7,
	output aout_8,
	output aout_9,
	output aout_10,
	output aout_11,
	output aout_12,
	output aout_13,
	output aout_14,
	output aout_15,
	output aout_16,
	output aout_17,
	output aout_18,
	output aout_19,
	output aout_20,
	output aout_21,
	output aout_22,
	output aout_23,
	output dsp16,
	output bigend,
	input sys_clk // Generated
);
wire d5_0;
wire d5_1;
wire d5_2;
wire d5_3;
wire d5_4;
wire d5_5;
wire d5_6;
wire d5_7;
wire d5_8;
wire d5_9;
wire d5_10;
wire d5_11;
wire d5_12;
wire d5_13;
wire d5_14;
wire d5_15;
wire d1_0;
wire d1_1;
wire d1_2;
wire d1_3;
wire d1_4;
wire d1_5;
wire d1_6;
wire d1_7;
wire d1_8;
wire d1_9;
wire d1_10;
wire d1_11;
wire d1_12;
wire d1_13;
wire d1_14;
wire d1_15;
wire d1_16;
wire d1_17;
wire d1_18;
wire d1_19;
wire d1_20;
wire d1_21;
wire d1_22;
wire d1_23;
wire d1_24;
wire d1_25;
wire d1_26;
wire d1_27;
wire d1_28;
wire d1_29;
wire d1_30;
wire d1_31;
wire d1a_8;
wire d1a_9;
wire d1a_10;
wire d1a_11;
wire d1a_12;
wire d1a_13;
wire d1a_14;
wire d1a_15;
wire d2_16;
wire d2_17;
wire d2_18;
wire d2_19;
wire d2_20;
wire d2_21;
wire d2_22;
wire d2_23;
wire d2_24;
wire d2_25;
wire d2_26;
wire d2_27;
wire d2_28;
wire d2_29;
wire d2_30;
wire d2_31;
wire d3_0;
wire d3_1;
wire d3_2;
wire d3_3;
wire d3_4;
wire d3_5;
wire d3_6;
wire d3_7;
wire d3_8;
wire d3_9;
wire d3_10;
wire d3_11;
wire d3_12;
wire d3_13;
wire d3_14;
wire d3_15;
wire d3_16;
wire d3_17;
wire d3_18;
wire d3_19;
wire d3_20;
wire d3_21;
wire d3_22;
wire d3_23;
wire d3_24;
wire d3_25;
wire d3_26;
wire d3_27;
wire d3_28;
wire d3_29;
wire d3_30;
wire d3_31;
wire d4_0;
wire d4_1;
wire d4_2;
wire d4_3;
wire d4_4;
wire d4_5;
wire d4_6;
wire d4_7;
wire d4_8;
wire d4_9;
wire d4_10;
wire d4_11;
wire d4_12;
wire d4_13;
wire d4_14;
wire d4_15;
wire d4a_0;
wire d4a_1;
wire d4a_2;
wire d4a_3;
wire d4a_4;
wire d4a_5;
wire d4a_6;
wire d4a_7;
wire d6_0;
wire d6_1;
wire d6_2;
wire d6_3;
wire d6_4;
wire d6_5;
wire d6_6;
wire d6_7;
wire d6_8;
wire d6_9;
wire d6_10;
wire d6_11;
wire d6_12;
wire d6_13;
wire d6_14;
wire d6_15;
wire ad_0;
wire ad_1;
wire ad_2;
wire ad_3;
wire ad_4;
wire ad_5;
wire ad_6;
wire ad_7;
wire ad_8;
wire ad_9;
wire ad_10;
wire ad_11;
wire ad_12;
wire ad_13;
wire ad_14;
wire ad_15;
wire ad_16;
wire ad_17;
wire ad_18;
wire ad_19;
wire ad_20;
wire ad_21;
wire ad_22;
wire ad_23;
wire as_1;
wire aouti_1;
wire aouti_14;

// JBUS.NET (44) - d5[0-15] : mx2
mx2 d5_from_0_to_15_inst_0
(
	.z /* OUT */ (d5_0),
	.a0 /* IN */ (din_0),
	.a1 /* IN */ (dr_0),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_1
(
	.z /* OUT */ (d5_1),
	.a0 /* IN */ (din_1),
	.a1 /* IN */ (dr_1),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_2
(
	.z /* OUT */ (d5_2),
	.a0 /* IN */ (din_2),
	.a1 /* IN */ (dr_2),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_3
(
	.z /* OUT */ (d5_3),
	.a0 /* IN */ (din_3),
	.a1 /* IN */ (dr_3),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_4
(
	.z /* OUT */ (d5_4),
	.a0 /* IN */ (din_4),
	.a1 /* IN */ (dr_4),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_5
(
	.z /* OUT */ (d5_5),
	.a0 /* IN */ (din_5),
	.a1 /* IN */ (dr_5),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_6
(
	.z /* OUT */ (d5_6),
	.a0 /* IN */ (din_6),
	.a1 /* IN */ (dr_6),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_7
(
	.z /* OUT */ (d5_7),
	.a0 /* IN */ (din_7),
	.a1 /* IN */ (dr_7),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_8
(
	.z /* OUT */ (d5_8),
	.a0 /* IN */ (din_8),
	.a1 /* IN */ (dr_8),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_9
(
	.z /* OUT */ (d5_9),
	.a0 /* IN */ (din_9),
	.a1 /* IN */ (dr_9),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_10
(
	.z /* OUT */ (d5_10),
	.a0 /* IN */ (din_10),
	.a1 /* IN */ (dr_10),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_11
(
	.z /* OUT */ (d5_11),
	.a0 /* IN */ (din_11),
	.a1 /* IN */ (dr_11),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_12
(
	.z /* OUT */ (d5_12),
	.a0 /* IN */ (din_12),
	.a1 /* IN */ (dr_12),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_13
(
	.z /* OUT */ (d5_13),
	.a0 /* IN */ (din_13),
	.a1 /* IN */ (dr_13),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_14
(
	.z /* OUT */ (d5_14),
	.a0 /* IN */ (din_14),
	.a1 /* IN */ (dr_14),
	.s /* IN */ (dren)
);
mx2 d5_from_0_to_15_inst_15
(
	.z /* OUT */ (d5_15),
	.a0 /* IN */ (din_15),
	.a1 /* IN */ (dr_15),
	.s /* IN */ (dren)
);

// JBUS.NET (48) - d1[0-31] : mx2
mx2 d1_from_0_to_31_inst_0
(
	.z /* OUT */ (d1_0),
	.a0 /* IN */ (wd_0),
	.a1 /* IN */ (din_0),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_1
(
	.z /* OUT */ (d1_1),
	.a0 /* IN */ (wd_1),
	.a1 /* IN */ (din_1),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_2
(
	.z /* OUT */ (d1_2),
	.a0 /* IN */ (wd_2),
	.a1 /* IN */ (din_2),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_3
(
	.z /* OUT */ (d1_3),
	.a0 /* IN */ (wd_3),
	.a1 /* IN */ (din_3),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_4
(
	.z /* OUT */ (d1_4),
	.a0 /* IN */ (wd_4),
	.a1 /* IN */ (din_4),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_5
(
	.z /* OUT */ (d1_5),
	.a0 /* IN */ (wd_5),
	.a1 /* IN */ (din_5),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_6
(
	.z /* OUT */ (d1_6),
	.a0 /* IN */ (wd_6),
	.a1 /* IN */ (din_6),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_7
(
	.z /* OUT */ (d1_7),
	.a0 /* IN */ (wd_7),
	.a1 /* IN */ (din_7),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_8
(
	.z /* OUT */ (d1_8),
	.a0 /* IN */ (wd_8),
	.a1 /* IN */ (din_8),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_9
(
	.z /* OUT */ (d1_9),
	.a0 /* IN */ (wd_9),
	.a1 /* IN */ (din_9),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_10
(
	.z /* OUT */ (d1_10),
	.a0 /* IN */ (wd_10),
	.a1 /* IN */ (din_10),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_11
(
	.z /* OUT */ (d1_11),
	.a0 /* IN */ (wd_11),
	.a1 /* IN */ (din_11),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_12
(
	.z /* OUT */ (d1_12),
	.a0 /* IN */ (wd_12),
	.a1 /* IN */ (din_12),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_13
(
	.z /* OUT */ (d1_13),
	.a0 /* IN */ (wd_13),
	.a1 /* IN */ (din_13),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_14
(
	.z /* OUT */ (d1_14),
	.a0 /* IN */ (wd_14),
	.a1 /* IN */ (din_14),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_15
(
	.z /* OUT */ (d1_15),
	.a0 /* IN */ (wd_15),
	.a1 /* IN */ (din_15),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_16
(
	.z /* OUT */ (d1_16),
	.a0 /* IN */ (wd_16),
	.a1 /* IN */ (din_16),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_17
(
	.z /* OUT */ (d1_17),
	.a0 /* IN */ (wd_17),
	.a1 /* IN */ (din_17),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_18
(
	.z /* OUT */ (d1_18),
	.a0 /* IN */ (wd_18),
	.a1 /* IN */ (din_18),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_19
(
	.z /* OUT */ (d1_19),
	.a0 /* IN */ (wd_19),
	.a1 /* IN */ (din_19),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_20
(
	.z /* OUT */ (d1_20),
	.a0 /* IN */ (wd_20),
	.a1 /* IN */ (din_20),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_21
(
	.z /* OUT */ (d1_21),
	.a0 /* IN */ (wd_21),
	.a1 /* IN */ (din_21),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_22
(
	.z /* OUT */ (d1_22),
	.a0 /* IN */ (wd_22),
	.a1 /* IN */ (din_22),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_23
(
	.z /* OUT */ (d1_23),
	.a0 /* IN */ (wd_23),
	.a1 /* IN */ (din_23),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_24
(
	.z /* OUT */ (d1_24),
	.a0 /* IN */ (wd_24),
	.a1 /* IN */ (din_24),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_25
(
	.z /* OUT */ (d1_25),
	.a0 /* IN */ (wd_25),
	.a1 /* IN */ (din_25),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_26
(
	.z /* OUT */ (d1_26),
	.a0 /* IN */ (wd_26),
	.a1 /* IN */ (din_26),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_27
(
	.z /* OUT */ (d1_27),
	.a0 /* IN */ (wd_27),
	.a1 /* IN */ (din_27),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_28
(
	.z /* OUT */ (d1_28),
	.a0 /* IN */ (wd_28),
	.a1 /* IN */ (din_28),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_29
(
	.z /* OUT */ (d1_29),
	.a0 /* IN */ (wd_29),
	.a1 /* IN */ (din_29),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_30
(
	.z /* OUT */ (d1_30),
	.a0 /* IN */ (wd_30),
	.a1 /* IN */ (din_30),
	.s /* IN */ (xdsrc)
);
mx2 d1_from_0_to_31_inst_31
(
	.z /* OUT */ (d1_31),
	.a0 /* IN */ (wd_31),
	.a1 /* IN */ (din_31),
	.s /* IN */ (xdsrc)
);

// JBUS.NET (52) - d1a[8-15] : mx2
mx2 d1a_from_8_to_15_inst_0
(
	.z /* OUT */ (d1a_8),
	.a0 /* IN */ (d1_8),
	.a1 /* IN */ (d1_0),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_1
(
	.z /* OUT */ (d1a_9),
	.a0 /* IN */ (d1_9),
	.a1 /* IN */ (d1_1),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_2
(
	.z /* OUT */ (d1a_10),
	.a0 /* IN */ (d1_10),
	.a1 /* IN */ (d1_2),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_3
(
	.z /* OUT */ (d1a_11),
	.a0 /* IN */ (d1_11),
	.a1 /* IN */ (d1_3),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_4
(
	.z /* OUT */ (d1a_12),
	.a0 /* IN */ (d1_12),
	.a1 /* IN */ (d1_4),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_5
(
	.z /* OUT */ (d1a_13),
	.a0 /* IN */ (d1_13),
	.a1 /* IN */ (d1_5),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_6
(
	.z /* OUT */ (d1a_14),
	.a0 /* IN */ (d1_14),
	.a1 /* IN */ (d1_6),
	.s /* IN */ (dmuxu_0)
);
mx2 d1a_from_8_to_15_inst_7
(
	.z /* OUT */ (d1a_15),
	.a0 /* IN */ (d1_15),
	.a1 /* IN */ (d1_7),
	.s /* IN */ (dmuxu_0)
);

// JBUS.NET (53) - d2[16-23] : mx2
mx2 d2_from_16_to_23_inst_0
(
	.z /* OUT */ (d2_16),
	.a0 /* IN */ (d1_16),
	.a1 /* IN */ (d1_0),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_1
(
	.z /* OUT */ (d2_17),
	.a0 /* IN */ (d1_17),
	.a1 /* IN */ (d1_1),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_2
(
	.z /* OUT */ (d2_18),
	.a0 /* IN */ (d1_18),
	.a1 /* IN */ (d1_2),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_3
(
	.z /* OUT */ (d2_19),
	.a0 /* IN */ (d1_19),
	.a1 /* IN */ (d1_3),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_4
(
	.z /* OUT */ (d2_20),
	.a0 /* IN */ (d1_20),
	.a1 /* IN */ (d1_4),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_5
(
	.z /* OUT */ (d2_21),
	.a0 /* IN */ (d1_21),
	.a1 /* IN */ (d1_5),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_6
(
	.z /* OUT */ (d2_22),
	.a0 /* IN */ (d1_22),
	.a1 /* IN */ (d1_6),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_16_to_23_inst_7
(
	.z /* OUT */ (d2_23),
	.a0 /* IN */ (d1_23),
	.a1 /* IN */ (d1_7),
	.s /* IN */ (dmuxu_1)
);

// JBUS.NET (54) - d2[24-31] : mx2
mx2 d2_from_24_to_31_inst_0
(
	.z /* OUT */ (d2_24),
	.a0 /* IN */ (d1_24),
	.a1 /* IN */ (d1a_8),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_1
(
	.z /* OUT */ (d2_25),
	.a0 /* IN */ (d1_25),
	.a1 /* IN */ (d1a_9),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_2
(
	.z /* OUT */ (d2_26),
	.a0 /* IN */ (d1_26),
	.a1 /* IN */ (d1a_10),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_3
(
	.z /* OUT */ (d2_27),
	.a0 /* IN */ (d1_27),
	.a1 /* IN */ (d1a_11),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_4
(
	.z /* OUT */ (d2_28),
	.a0 /* IN */ (d1_28),
	.a1 /* IN */ (d1a_12),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_5
(
	.z /* OUT */ (d2_29),
	.a0 /* IN */ (d1_29),
	.a1 /* IN */ (d1a_13),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_6
(
	.z /* OUT */ (d2_30),
	.a0 /* IN */ (d1_30),
	.a1 /* IN */ (d1a_14),
	.s /* IN */ (dmuxu_1)
);
mx2 d2_from_24_to_31_inst_7
(
	.z /* OUT */ (d2_31),
	.a0 /* IN */ (d1_31),
	.a1 /* IN */ (d1a_15),
	.s /* IN */ (dmuxu_1)
);

// JBUS.NET (58) - d3[0-7] : stlatch
stlatch d3_from_0_to_7_inst_0
(
	.d1 /* OUT */ (d3_0),
	.d /* IN */ (d1_0),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_1
(
	.d1 /* OUT */ (d3_1),
	.d /* IN */ (d1_1),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_2
(
	.d1 /* OUT */ (d3_2),
	.d /* IN */ (d1_2),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_3
(
	.d1 /* OUT */ (d3_3),
	.d /* IN */ (d1_3),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_4
(
	.d1 /* OUT */ (d3_4),
	.d /* IN */ (d1_4),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_5
(
	.d1 /* OUT */ (d3_5),
	.d /* IN */ (d1_5),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_6
(
	.d1 /* OUT */ (d3_6),
	.d /* IN */ (d1_6),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_0_to_7_inst_7
(
	.d1 /* OUT */ (d3_7),
	.d /* IN */ (d1_7),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);

// JBUS.NET (59) - d3[8-15] : stlatch
stlatch d3_from_8_to_15_inst_0
(
	.d1 /* OUT */ (d3_8),
	.d /* IN */ (d1a_8),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_1
(
	.d1 /* OUT */ (d3_9),
	.d /* IN */ (d1a_9),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_2
(
	.d1 /* OUT */ (d3_10),
	.d /* IN */ (d1a_10),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_3
(
	.d1 /* OUT */ (d3_11),
	.d /* IN */ (d1a_11),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_4
(
	.d1 /* OUT */ (d3_12),
	.d /* IN */ (d1a_12),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_5
(
	.d1 /* OUT */ (d3_13),
	.d /* IN */ (d1a_13),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_6
(
	.d1 /* OUT */ (d3_14),
	.d /* IN */ (d1a_14),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_8_to_15_inst_7
(
	.d1 /* OUT */ (d3_15),
	.d /* IN */ (d1a_15),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_0),
	.sys_clk(sys_clk) // Generated
);

// JBUS.NET (60) - d3[16-31] : stlatch
stlatch d3_from_16_to_31_inst_0
(
	.d1 /* OUT */ (d3_16),
	.d /* IN */ (d2_16),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_1
(
	.d1 /* OUT */ (d3_17),
	.d /* IN */ (d2_17),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_2
(
	.d1 /* OUT */ (d3_18),
	.d /* IN */ (d2_18),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_3
(
	.d1 /* OUT */ (d3_19),
	.d /* IN */ (d2_19),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_4
(
	.d1 /* OUT */ (d3_20),
	.d /* IN */ (d2_20),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_5
(
	.d1 /* OUT */ (d3_21),
	.d /* IN */ (d2_21),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_6
(
	.d1 /* OUT */ (d3_22),
	.d /* IN */ (d2_22),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_7
(
	.d1 /* OUT */ (d3_23),
	.d /* IN */ (d2_23),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_8
(
	.d1 /* OUT */ (d3_24),
	.d /* IN */ (d2_24),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_9
(
	.d1 /* OUT */ (d3_25),
	.d /* IN */ (d2_25),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_10
(
	.d1 /* OUT */ (d3_26),
	.d /* IN */ (d2_26),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_11
(
	.d1 /* OUT */ (d3_27),
	.d /* IN */ (d2_27),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_12
(
	.d1 /* OUT */ (d3_28),
	.d /* IN */ (d2_28),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_13
(
	.d1 /* OUT */ (d3_29),
	.d /* IN */ (d2_29),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_14
(
	.d1 /* OUT */ (d3_30),
	.d /* IN */ (d2_30),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);
stlatch d3_from_16_to_31_inst_15
(
	.d1 /* OUT */ (d3_31),
	.d /* IN */ (d2_31),
	.clk /* IN */ (clk),
	.en /* IN */ (dinlatch_1),
	.sys_clk(sys_clk) // Generated
);

// JBUS.NET (64) - d4[0-15] : mx2
mx2 d4_from_0_to_15_inst_0
(
	.z /* OUT */ (d4_0),
	.a0 /* IN */ (d3_0),
	.a1 /* IN */ (d3_16),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_1
(
	.z /* OUT */ (d4_1),
	.a0 /* IN */ (d3_1),
	.a1 /* IN */ (d3_17),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_2
(
	.z /* OUT */ (d4_2),
	.a0 /* IN */ (d3_2),
	.a1 /* IN */ (d3_18),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_3
(
	.z /* OUT */ (d4_3),
	.a0 /* IN */ (d3_3),
	.a1 /* IN */ (d3_19),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_4
(
	.z /* OUT */ (d4_4),
	.a0 /* IN */ (d3_4),
	.a1 /* IN */ (d3_20),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_5
(
	.z /* OUT */ (d4_5),
	.a0 /* IN */ (d3_5),
	.a1 /* IN */ (d3_21),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_6
(
	.z /* OUT */ (d4_6),
	.a0 /* IN */ (d3_6),
	.a1 /* IN */ (d3_22),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_7
(
	.z /* OUT */ (d4_7),
	.a0 /* IN */ (d3_7),
	.a1 /* IN */ (d3_23),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_8
(
	.z /* OUT */ (d4_8),
	.a0 /* IN */ (d3_8),
	.a1 /* IN */ (d3_24),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_9
(
	.z /* OUT */ (d4_9),
	.a0 /* IN */ (d3_9),
	.a1 /* IN */ (d3_25),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_10
(
	.z /* OUT */ (d4_10),
	.a0 /* IN */ (d3_10),
	.a1 /* IN */ (d3_26),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_11
(
	.z /* OUT */ (d4_11),
	.a0 /* IN */ (d3_11),
	.a1 /* IN */ (d3_27),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_12
(
	.z /* OUT */ (d4_12),
	.a0 /* IN */ (d3_12),
	.a1 /* IN */ (d3_28),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_13
(
	.z /* OUT */ (d4_13),
	.a0 /* IN */ (d3_13),
	.a1 /* IN */ (d3_29),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_14
(
	.z /* OUT */ (d4_14),
	.a0 /* IN */ (d3_14),
	.a1 /* IN */ (d3_30),
	.s /* IN */ (dmuxd_1)
);
mx2 d4_from_0_to_15_inst_15
(
	.z /* OUT */ (d4_15),
	.a0 /* IN */ (d3_15),
	.a1 /* IN */ (d3_31),
	.s /* IN */ (dmuxd_1)
);

// JBUS.NET (65) - d4a[0-7] : mx2
mx2 d4a_from_0_to_7_inst_0
(
	.z /* OUT */ (d4a_0),
	.a0 /* IN */ (d4_0),
	.a1 /* IN */ (d4_8),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_1
(
	.z /* OUT */ (d4a_1),
	.a0 /* IN */ (d4_1),
	.a1 /* IN */ (d4_9),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_2
(
	.z /* OUT */ (d4a_2),
	.a0 /* IN */ (d4_2),
	.a1 /* IN */ (d4_10),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_3
(
	.z /* OUT */ (d4a_3),
	.a0 /* IN */ (d4_3),
	.a1 /* IN */ (d4_11),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_4
(
	.z /* OUT */ (d4a_4),
	.a0 /* IN */ (d4_4),
	.a1 /* IN */ (d4_12),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_5
(
	.z /* OUT */ (d4a_5),
	.a0 /* IN */ (d4_5),
	.a1 /* IN */ (d4_13),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_6
(
	.z /* OUT */ (d4a_6),
	.a0 /* IN */ (d4_6),
	.a1 /* IN */ (d4_14),
	.s /* IN */ (dmuxd_0)
);
mx2 d4a_from_0_to_7_inst_7
(
	.z /* OUT */ (d4a_7),
	.a0 /* IN */ (d4_7),
	.a1 /* IN */ (d4_15),
	.s /* IN */ (dmuxd_0)
);

// JBUS.NET (69) - d6[0-7] : mx2
mx2 d6_from_0_to_7_inst_0
(
	.z /* OUT */ (d6_0),
	.a0 /* IN */ (d5_0),
	.a1 /* IN */ (d4a_0),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_1
(
	.z /* OUT */ (d6_1),
	.a0 /* IN */ (d5_1),
	.a1 /* IN */ (d4a_1),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_2
(
	.z /* OUT */ (d6_2),
	.a0 /* IN */ (d5_2),
	.a1 /* IN */ (d4a_2),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_3
(
	.z /* OUT */ (d6_3),
	.a0 /* IN */ (d5_3),
	.a1 /* IN */ (d4a_3),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_4
(
	.z /* OUT */ (d6_4),
	.a0 /* IN */ (d5_4),
	.a1 /* IN */ (d4a_4),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_5
(
	.z /* OUT */ (d6_5),
	.a0 /* IN */ (d5_5),
	.a1 /* IN */ (d4a_5),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_6
(
	.z /* OUT */ (d6_6),
	.a0 /* IN */ (d5_6),
	.a1 /* IN */ (d4a_6),
	.s /* IN */ (masterdata)
);
mx2 d6_from_0_to_7_inst_7
(
	.z /* OUT */ (d6_7),
	.a0 /* IN */ (d5_7),
	.a1 /* IN */ (d4a_7),
	.s /* IN */ (masterdata)
);

// JBUS.NET (70) - d6[8-15] : mx2
mx2 d6_from_8_to_15_inst_0
(
	.z /* OUT */ (d6_8),
	.a0 /* IN */ (d5_8),
	.a1 /* IN */ (d4_8),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_1
(
	.z /* OUT */ (d6_9),
	.a0 /* IN */ (d5_9),
	.a1 /* IN */ (d4_9),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_2
(
	.z /* OUT */ (d6_10),
	.a0 /* IN */ (d5_10),
	.a1 /* IN */ (d4_10),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_3
(
	.z /* OUT */ (d6_11),
	.a0 /* IN */ (d5_11),
	.a1 /* IN */ (d4_11),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_4
(
	.z /* OUT */ (d6_12),
	.a0 /* IN */ (d5_12),
	.a1 /* IN */ (d4_12),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_5
(
	.z /* OUT */ (d6_13),
	.a0 /* IN */ (d5_13),
	.a1 /* IN */ (d4_13),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_6
(
	.z /* OUT */ (d6_14),
	.a0 /* IN */ (d5_14),
	.a1 /* IN */ (d4_14),
	.s /* IN */ (masterdata)
);
mx2 d6_from_8_to_15_inst_7
(
	.z /* OUT */ (d6_15),
	.a0 /* IN */ (d5_15),
	.a1 /* IN */ (d4_15),
	.s /* IN */ (masterdata)
);

// JBUS.NET (74) - dout[0-15] : nivh
assign dout_0 = d6_0;
assign dout_1 = d6_1;
assign dout_2 = d6_2;
assign dout_3 = d6_3;
assign dout_4 = d6_4;
assign dout_5 = d6_5;
assign dout_6 = d6_6;
assign dout_7 = d6_7;
assign dout_8 = d6_8;
assign dout_9 = d6_9;
assign dout_10 = d6_10;
assign dout_11 = d6_11;
assign dout_12 = d6_12;
assign dout_13 = d6_13;
assign dout_14 = d6_14;
assign dout_15 = d6_15;

// JBUS.NET (75) - dout[16-31] : nivm
assign dout_16 = d3_16;
assign dout_17 = d3_17;
assign dout_18 = d3_18;
assign dout_19 = d3_19;
assign dout_20 = d3_20;
assign dout_21 = d3_21;
assign dout_22 = d3_22;
assign dout_23 = d3_23;
assign dout_24 = d3_24;
assign dout_25 = d3_25;
assign dout_26 = d3_26;
assign dout_27 = d3_27;
assign dout_28 = d3_28;
assign dout_29 = d3_29;
assign dout_30 = d3_30;
assign dout_31 = d3_31;

// JBUS.NET (79) - dsp16 : ldp1q
ldp1q dsp16_inst
(
	.q /* OUT */ (dsp16),
	.d /* IN */ (cfg_0),
	.g /* IN */ (cfgw),
	.sys_clk(sys_clk) // Generated
);

// JBUS.NET (80) - bigend : ldp1q
ldp1q bigend_inst
(
	.q /* OUT */ (bigend),
	.d /* IN */ (cfg_1),
	.g /* IN */ (cfgw),
	.sys_clk(sys_clk) // Generated
);

// JBUS.NET (86) - ad[0-23] : slatch
j_slatch ad_from_0_to_23_inst_0
(
	.q /* OUT */ (ad_0),
	.d /* IN */ (a_0),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_1
(
	.q /* OUT */ (ad_1),
	.d /* IN */ (a_1),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_2
(
	.q /* OUT */ (ad_2),
	.d /* IN */ (a_2),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_3
(
	.q /* OUT */ (ad_3),
	.d /* IN */ (a_3),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_4
(
	.q /* OUT */ (ad_4),
	.d /* IN */ (a_4),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_5
(
	.q /* OUT */ (ad_5),
	.d /* IN */ (a_5),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_6
(
	.q /* OUT */ (ad_6),
	.d /* IN */ (a_6),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_7
(
	.q /* OUT */ (ad_7),
	.d /* IN */ (a_7),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_8
(
	.q /* OUT */ (ad_8),
	.d /* IN */ (a_8),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_9
(
	.q /* OUT */ (ad_9),
	.d /* IN */ (a_9),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_10
(
	.q /* OUT */ (ad_10),
	.d /* IN */ (a_10),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_11
(
	.q /* OUT */ (ad_11),
	.d /* IN */ (a_11),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_12
(
	.q /* OUT */ (ad_12),
	.d /* IN */ (a_12),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_13
(
	.q /* OUT */ (ad_13),
	.d /* IN */ (a_13),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_14
(
	.q /* OUT */ (ad_14),
	.d /* IN */ (a_14),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_15
(
	.q /* OUT */ (ad_15),
	.d /* IN */ (a_15),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_16
(
	.q /* OUT */ (ad_16),
	.d /* IN */ (a_16),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_17
(
	.q /* OUT */ (ad_17),
	.d /* IN */ (a_17),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_18
(
	.q /* OUT */ (ad_18),
	.d /* IN */ (a_18),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_19
(
	.q /* OUT */ (ad_19),
	.d /* IN */ (a_19),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_20
(
	.q /* OUT */ (ad_20),
	.d /* IN */ (a_20),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_21
(
	.q /* OUT */ (ad_21),
	.d /* IN */ (a_21),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_22
(
	.q /* OUT */ (ad_22),
	.d /* IN */ (a_22),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);
j_slatch ad_from_0_to_23_inst_23
(
	.q /* OUT */ (ad_23),
	.d /* IN */ (a_23),
	.clk /* IN */ (clk),
	.en /* IN */ (ack),
	.sys_clk(sys_clk) // Generated
);

// JBUS.NET (88) - as[1] : or2
assign as_1 = ad_1 | seta1;

// JBUS.NET (90) - aout[0] : mx2
mx2 aout_index_0_inst
(
	.z /* OUT */ (aout_0),
	.a0 /* IN */ (ad_0),
	.a1 /* IN */ (ain_0),
	.s /* IN */ (ainen)
);

// JBUS.NET (91) - aouti[1] : mx2
mx2 aouti_index_1_inst
(
	.z /* OUT */ (aouti_1),
	.a0 /* IN */ (as_1),
	.a1 /* IN */ (ain_1),
	.s /* IN */ (ainen)
);

// JBUS.NET (92) - aout[1] : nivu
assign aout_1 = aouti_1;

// JBUS.NET (93) - aout[2-13] : mx2
mx2 aout_from_2_to_13_inst_0
(
	.z /* OUT */ (aout_2),
	.a0 /* IN */ (ad_2),
	.a1 /* IN */ (ain_2),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_1
(
	.z /* OUT */ (aout_3),
	.a0 /* IN */ (ad_3),
	.a1 /* IN */ (ain_3),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_2
(
	.z /* OUT */ (aout_4),
	.a0 /* IN */ (ad_4),
	.a1 /* IN */ (ain_4),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_3
(
	.z /* OUT */ (aout_5),
	.a0 /* IN */ (ad_5),
	.a1 /* IN */ (ain_5),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_4
(
	.z /* OUT */ (aout_6),
	.a0 /* IN */ (ad_6),
	.a1 /* IN */ (ain_6),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_5
(
	.z /* OUT */ (aout_7),
	.a0 /* IN */ (ad_7),
	.a1 /* IN */ (ain_7),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_6
(
	.z /* OUT */ (aout_8),
	.a0 /* IN */ (ad_8),
	.a1 /* IN */ (ain_8),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_7
(
	.z /* OUT */ (aout_9),
	.a0 /* IN */ (ad_9),
	.a1 /* IN */ (ain_9),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_8
(
	.z /* OUT */ (aout_10),
	.a0 /* IN */ (ad_10),
	.a1 /* IN */ (ain_10),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_9
(
	.z /* OUT */ (aout_11),
	.a0 /* IN */ (ad_11),
	.a1 /* IN */ (ain_11),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_10
(
	.z /* OUT */ (aout_12),
	.a0 /* IN */ (ad_12),
	.a1 /* IN */ (ain_12),
	.s /* IN */ (ainen)
);
mx2 aout_from_2_to_13_inst_11
(
	.z /* OUT */ (aout_13),
	.a0 /* IN */ (ad_13),
	.a1 /* IN */ (ain_13),
	.s /* IN */ (ainen)
);

// JBUS.NET (94) - aouti[14] : mx2
mx2 aouti_index_14_inst
(
	.z /* OUT */ (aouti_14),
	.a0 /* IN */ (ad_14),
	.a1 /* IN */ (ain_14),
	.s /* IN */ (ainen)
);

// JBUS.NET (95) - aout[14] : nivh
assign aout_14 = aouti_14;

// JBUS.NET (96) - aout[15-23] : mx2
mx2 aout_from_15_to_23_inst_0
(
	.z /* OUT */ (aout_15),
	.a0 /* IN */ (ad_15),
	.a1 /* IN */ (ain_15),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_1
(
	.z /* OUT */ (aout_16),
	.a0 /* IN */ (ad_16),
	.a1 /* IN */ (ain_16),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_2
(
	.z /* OUT */ (aout_17),
	.a0 /* IN */ (ad_17),
	.a1 /* IN */ (ain_17),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_3
(
	.z /* OUT */ (aout_18),
	.a0 /* IN */ (ad_18),
	.a1 /* IN */ (ain_18),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_4
(
	.z /* OUT */ (aout_19),
	.a0 /* IN */ (ad_19),
	.a1 /* IN */ (ain_19),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_5
(
	.z /* OUT */ (aout_20),
	.a0 /* IN */ (ad_20),
	.a1 /* IN */ (ain_20),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_6
(
	.z /* OUT */ (aout_21),
	.a0 /* IN */ (ad_21),
	.a1 /* IN */ (ain_21),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_7
(
	.z /* OUT */ (aout_22),
	.a0 /* IN */ (ad_22),
	.a1 /* IN */ (ain_22),
	.s /* IN */ (ainen)
);
mx2 aout_from_15_to_23_inst_8
(
	.z /* OUT */ (aout_23),
	.a0 /* IN */ (ad_23),
	.a1 /* IN */ (ain_23),
	.s /* IN */ (ainen)
);
endmodule
/* verilator lint_on LITENDIAN */
