module pll50 (
	input inclk0,
	output c0,
	output c1,
	output c2,
	output c3);

assign c0 = inclk0;
assign c1 = inclk0;
assign c2 = inclk0;
assign c3 = inclk0;

endmodule

